library verilog;
use verilog.vl_types.all;
entity controller is
    generic(
        state_reset     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        read            : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        decode          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        adi_execute     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        regw_frm_aluout : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        i_type_load     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        lhi_execute     : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        i_type_store    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        branch_compare  : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        br_check        : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        br_yes          : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        jmp_add         : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        jmp_store_pc    : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        add             : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        nanda           : vl_logic_vector(0 to 15) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        jlr             : vl_logic_vector(0 to 15) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        lw_execute      : vl_logic_vector(0 to 15) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        sw_execute      : vl_logic_vector(0 to 15) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        LM1             : vl_logic_vector(0 to 15) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        LM2             : vl_logic_vector(0 to 15) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        LM3             : vl_logic_vector(0 to 15) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        SM              : vl_logic_vector(0 to 15) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0)
    );
    port(
        reset           : in     vl_logic;
        clk             : in     vl_logic;
        mem_read        : out    vl_logic;
        mem_write       : out    vl_logic;
        R_pc            : out    vl_logic_vector(1 downto 0);
        alusrc_a        : out    vl_logic;
        alusrc_b        : out    vl_logic_vector(1 downto 0);
        regdst          : out    vl_logic_vector(1 downto 0);
        reg_w           : out    vl_logic;
        b_c             : out    vl_logic_vector(1 downto 0);
        memtoreg        : out    vl_logic_vector(1 downto 0);
        i_d             : out    vl_logic;
        ir_w            : out    vl_logic;
        alu_op          : out    vl_logic_vector(1 downto 0);
        inst            : in     vl_logic_vector(15 downto 0);
        car_zer         : in     vl_logic_vector(1 downto 0);
        st              : out    vl_logic_vector(15 downto 0);
        ccr_update      : out    vl_logic;
        enbl            : out    vl_logic;
        count           : in     vl_logic_vector(2 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of state_reset : constant is 1;
    attribute mti_svvh_generic_type of read : constant is 1;
    attribute mti_svvh_generic_type of decode : constant is 1;
    attribute mti_svvh_generic_type of adi_execute : constant is 1;
    attribute mti_svvh_generic_type of regw_frm_aluout : constant is 1;
    attribute mti_svvh_generic_type of i_type_load : constant is 1;
    attribute mti_svvh_generic_type of lhi_execute : constant is 1;
    attribute mti_svvh_generic_type of i_type_store : constant is 1;
    attribute mti_svvh_generic_type of branch_compare : constant is 1;
    attribute mti_svvh_generic_type of br_check : constant is 1;
    attribute mti_svvh_generic_type of br_yes : constant is 1;
    attribute mti_svvh_generic_type of jmp_add : constant is 1;
    attribute mti_svvh_generic_type of jmp_store_pc : constant is 1;
    attribute mti_svvh_generic_type of add : constant is 1;
    attribute mti_svvh_generic_type of nanda : constant is 1;
    attribute mti_svvh_generic_type of jlr : constant is 1;
    attribute mti_svvh_generic_type of lw_execute : constant is 1;
    attribute mti_svvh_generic_type of sw_execute : constant is 1;
    attribute mti_svvh_generic_type of LM1 : constant is 1;
    attribute mti_svvh_generic_type of LM2 : constant is 1;
    attribute mti_svvh_generic_type of LM3 : constant is 1;
    attribute mti_svvh_generic_type of SM : constant is 1;
end controller;
