module memory(clk, address, wrdata, dataout, mem_write, mem_read);
input [15:0]address;
input [15:0]wrdata;
input clk;
input  mem_read;
input  mem_write;
output reg[15:0] dataout;
reg [15:0] mem[63:0];	





initial begin
mem[0] =16'b1000000000011100;
mem[1] =16'b0100100110000101;
mem[2] =16'b0001000110111101;
mem[3] =16'b0100110110000101;
mem[4] =16'b0110000000000011;
mem[5] =16'b0001010000000000;
mem[6] =16'b0010000001011000;
mem[7] =16'b0010011011011000;
mem[8] =16'b0001011011000000;
mem[9] =16'b0000100010100001;
mem[10] =16'b0000000000000000;
mem[11] =16'b0010110110110010;
mem[12] =16'b1100110101111001;
mem[13] =16'b0101100101010110;

mem[20] =16'b0000000000000001;
mem[21] =16'b0000000000101111;
mem[22] =16'b0000000000000000;
mem[23] =16'b0000000000000101;
mem[24] =16'b0000000000000010;


mem[29] =16'b0001011011000001;
mem[30] =16'b0001110110010111;
mem[31] =16'b0101000110000100;
mem[32] =16'b0100000110000000;
mem[33] =16'b0100001110000001;
mem[34] =16'b1100101001001011;
mem[35] =16'b0000000010010000;
mem[36] =16'b0000011100100010;
mem[37] =16'b0001001001111111;
mem[38] =16'b0001111111111011;


mem[46] =16'b0001000110000010;
mem[47] =16'b0111000000010100;
mem[48] =16'b0001011011111111;
mem[49] =16'b0101011110000101;
mem[50] =16'b0100111110000100;
end
//initial begin
//mem[0] =16'b1000001000000001;
//mem[1] =16'b0100100110000101;
//mem[2] =16'b0100110110000101;
//mem[3] =16'b0100000101010100;//beq
//mem[4] =16'b0100001101010101;//add
//mem[5] =16'b1100101001000011;//beq
//mem[6] =16'b0010000000000100;
//mem[7] =16'b0010000111100100;
//mem[8] =16'b1100101001000010;
//mem[9] =16'b0010000000000100;
//mem[10] =16'b0010000000000100;
//mem[11] =16'b0010000000000100;
//mem[12] =16'b0010000000000100;
//mem[13] =16'b0111000001000110;
//mem[14] =16'b0010000000000100;
//mem[15] =16'b0010000000000100;
//end

//assign dataout=(mem_read==1'b1)?mem[address]:16'h0000;

always @(*) begin
	
	if(mem_read==1'b1)
		begin dataout = mem[address]; end
	else dataout = 16'b0;
end	
	

	
always @(posedge clk) begin
	
	if(mem_write==1'b1)
		begin mem[address] = wrdata; end
	

end
endmodule










